// SPDX-FileCopyrightText: (c) 2024  Parallel Architectures Group (GAP) <carherlu@upv.edu.es>
// SPDX-License-Identifier: MIT
//
//
// @file single_unit_network_interface_test_pkg.sv 
// @author Rafael Tornero (ratorga@disca.upv.es)
// @date March 05th, 2024
//
// @title Single Unit Network Interface test package
//
package single_unit_network_interface_test_pkg;
  
  import single_unit_network_interface_env_pkg::*;
  
endpackage
