`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////
// (c) Copyright 2012 - 2017  Parallel Architectures Group (GAP)
// Department of Computing Engineering (DISCA)
// Universitat Politecnica de Valencia (UPV)
// Valencia, Spain
// All rights reserved.
// 
// All code contained herein is, and remains the property of
// Parallel Architectures Group. The intellectual and technical concepts
// contained herein are proprietary to Parallel Architectures Group and 
// are protected by trade secret or copyright law.
// Dissemination of this code or reproduction of this material is 
// strictly forbidden unless prior written permission is obtained
// from Parallel Architectures Group.
//
// THIS SOFTWARE IS MADE AVAILABLE "AS IS" AND IT IS NOT INTENDED FOR USE
// IN WHICH THE FAILURE OF THE SOFTWARE COULD LEAD TO DEATH, PERSONAL INJURY,
// OR SEVERE PHYSICAL OR ENVIRONMENTAL DAMAGE.
// 
// contact: jflich@disca.upv.es
//-----------------------------------------------------------------------------
//
// Company:  GAP (UPV)  
// Engineer: T. Piconell (tompic@gap.upv.es)
// 
// Create Date: 
// Design Name: 
// Module Name: 
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//
//  
//
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////

// This module implements a fixed n-bit priority arbiter where the number of bits can be specified as a parameter (NUM_ARBITER_PORTS)
module FPA #(
  parameter NUM_ARBITER_PORTS = 1  // number of arbiter ports
)(
  input  [NUM_ARBITER_PORTS-1 : 0] vector_in,  // input vector (token requests)
  output [NUM_ARBITER_PORTS-1 : 0] vector_out  // output vector (grants)
);

  genvar j;
  generate
    assign vector_out[0] = vector_in[0];
    for( j=1; j<NUM_ARBITER_PORTS;j = j+1) begin : LOOP
        assign vector_out[j] = (vector_in[j]) & (~|vector_in[(j-1):0]);
    end
 endgenerate
endmodule
